/**********************************************
 Author: Rohit Srinivas R G, M Kapil Shyam
 Email: CS23Z002@smail.iitm.ac.in, CS23Z064@smail.iitm.ac.in
**********************************************/

package Testbench;

// ================================================================
// Project imports


// ================================================================

interface Ifc_Testbench;
  
endinterface

(* synthesize *)
module mkTestbench (Ifc_Testbench);

   
endmodule

// ================================================================

endpackage
           
